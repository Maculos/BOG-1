/*
RV64I CPU Project
Module is based on version 20191213 of the Unprivileged RISC-V ISA Chapter(s) 
XLEN = 64;
*/

`ifndef regfile
`define regfile

module regfile (
    input clock,
);





endmodule

`endif